BZh91AY&SY(VMN B߀Py��g߰����Px= fd
 e���z@�  � 4hɉ�	���0 �`�0�! ��$z�5O&�M�� �z��2b`b0#L1&L0H����&SFҙ1=MA��M���$(E�#"�z������?�
Ͱp
A��쳂�d �hX`z�F��:��۰
~&ӌmN�#�����Ni��7�K(�Ƴ��J���ii{�2�yz�G=�ݞV0��i�H�w���q<ͱ�Aa��"$�:"!#�����J�e &41�<���d.?MS��V.2гT��1[g���.:܀�+�^V5��:q����.2�����\�Y�ة[�mNQa��������{k��6zث�eT��!�n��[������vl`�X���5�����^׍�y��f�4��M6z�g
ao(w�������C@���܎� �i�U��]d�S�ܧW9��Y�+0�d	T
:�m%ͨ�G��DF���7�l���S%r�q��r.�����f�����X'G���.8A����Rf)��-� ��B���l`/�A�9ȇ*v���s��E�=�����_�u��H3����Љ6��8]|�=y;�NĽ�i�Go[���2��i�j;��u�g$��n!vG��_�qQYHù4�� p52L�)Z���,3UJ�% ����K�^�B�Ƣ[�&z�a��5��1H�>}y�M�M�\:rE_�F��@U^��_ۖ�̑�I����@]*\ǈ-�'#<!q5Xq����6"�)q��w���&�) cD＂=vW������:B+x���ăTɈPR�A�	�~ .b"6�+,"û}"�u�Dg����� �����AmKD�)C�hcFތ�W�Q0�4q�E(�e(�ഈ[��1Dن�jT�
k,5OM2(	��� �y���r��-k&,��O1�̒w�"�mC�PU���	�RdA*��󍍅�*>�lF����)�B�jp